`default_nettype none
`timescale 1ms / 10ns

module logicelement_tb;

  localparam int LUT_SIZE = 16;
  localparam int SEL_WIDTH = $clog2(LUT_SIZE);

  // Inputs
  logic clk, en, nrst;
  logic le_clk, le_en, le_nrst;
  logic [SEL_WIDTH-1:0] select;
  logic config_data_in, config_en, config_data_out; // +1 for mode
  int test_case;

  // Output
  logic le_out;

  // DUT
  logicelement #(.LUT_SIZE(LUT_SIZE)) dut (
    .clk(clk),
    .en(en),
    .nrst(nrst),
    .le_clk(le_clk),
    .le_en(le_en),
    .le_nrst(le_nrst),
    .select(select),
    .config_data_in(config_data_in),
    .config_en(config_en),
    .config_data_out(config_data_out),
    .le_out(le_out)
  );

  // Clock generation
  initial le_clk = 0;
  always #2 le_clk = ~le_clk; // 10ns clock period

  task le_reset();
    begin
      le_nrst = 0; le_en = 1; select = 0;
      #1;
      le_nrst = 1;
      #1;
    end
  endtask

  task reset();
    begin
      nrst = 0; en = 1; config_en = 0; config_data_in = 0; clk = 0;
      #1;
      nrst = 1;
      config_en = 1;
      #1;
    end
  endtask

  task cram(logic [(LUT_SIZE + 1) - 1:0] data);
    begin
      config_en = 1; //allow configuration
      for (int i = LUT_SIZE + 1; i > 0; i --) begin
        clk = 0;
        config_data_in = data[i - 1]; //MSB first
        #1;
        clk = 1;
        #1;
      end
      config_en = 0;
      le_reset();
    end
  endtask

  // LUT: Implement function: f(select) = select[0] ^ select[1] (for example)
  function automatic [LUT_SIZE-1:0] make_xor_lut();
    int i;
    logic [LUT_SIZE-1:0] lut;
    begin
      for (i = 0; i < LUT_SIZE; i++) begin
        lut[i] = ^i; // XOR of lower 2 bits of select
      end
      return lut;
    end
  endfunction

  logic [LUT_SIZE-1:0] xor_lut = make_xor_lut();

  initial begin

    $dumpfile("waves/logicelement.vcd"); //change the vcd vile name to your source file name
    $dumpvars(0, logicelement_tb);

    $display("Starting testbench...");
    le_reset();
    reset();
    test_case = 0;

    // === Test 1: Combinational Mode ===
    $display("Test 1: Combinational mode");
    test_case = 1;
    cram ({1'b0, xor_lut});
    for (int i = 0; i < LUT_SIZE; i++) begin
      select = i;
      #1; // allow propagation
      assert (le_out == xor_lut[i]) else
        $error("FAIL: select=%0d, expected=%0b, got=%0b", i, xor_lut[i], le_out);
    end

    le_reset();
    reset();

    // === Test 2: Registered Mode ===
    $display("Test 2: Registered (DFF) mode");
    test_case = 2;
    cram({1'b1, xor_lut});

    for (int i = 0; i < LUT_SIZE; i++) begin
      select = i;
      #2;
    end

    le_reset();
    reset();

    // === Test 3: DFF Hold Behavior ===
    $display("Test 3: Registered mode, en=0 (hold)");
    test_case = 3;
    cram({1'b1, 16'd1});
    #2
    select = 0;
    #1
    le_en = 0;
    #1
    select = select + 1; // change select, but en=0
    #10
    assert (le_out == 1) else
      $error("FAIL: DFF should hold value when en=0");

    $display("All tests completed.");
    $finish;
  end

endmodule
